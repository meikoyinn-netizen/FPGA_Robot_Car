`timescale 1ns / 1ps

module tb_my_pc_reg;

    // ==========================================
    // 1. 定义信号
    // ==========================================
    // 输入信号 (用 reg，因为要在 initial 块里赋值)
    reg clk;
    reg rst_n;
    reg stall;
    reg jump_flag;
    reg [31:0] jump_addr;

    // 输出信号 (用 wire，因为是连接模块的输出)
    wire [31:0] pc;

    // ==========================================
    // 2. 实例化被测模块 (把你的 PC 接上去)
    // ==========================================
    my_pc_reg uut (
        .clk(clk),
        .rst_n(rst_n),
        .stall(stall),
        .jump_flag(jump_flag),
        .jump_addr(jump_addr),
        .pc(pc)
    );

    // ==========================================
    // 3. 产生时钟 (模拟 50MHz 晶振)
    // ==========================================
    initial begin
        clk = 0;
        // 每 10ns 翻转一次，周期 20ns
        forever #10 clk = ~clk; 
    end

    // ==========================================
    // 4. 测试剧本
    // ==========================================
    initial begin
        // --- 初始化状态 ---
        rst_n = 0;      // 按下复位键
        stall = 0;
        jump_flag = 0;
        jump_addr = 0;

        // 等待 100ns，看看 PC 是不是归零了
        #100;
        
        // --- 场景 1: 正常计数 ---
        rst_n = 1;      // 松开复位，PC 应该开始跑 (0, 4, 8, 12...)
        #100;           // 让它跑 5 个周期

        // --- 场景 2: 测试暂停 (Stall) ---
        stall = 1;      // 喊停！PC 应该保持不动
        #60;            // 停一会儿
        stall = 0;      // 继续跑
        #60;

        // --- 场景 3: 测试跳转 (Jump) ---
        jump_addr = 32'h8000_1000; // 设定目标地址
        jump_flag = 1;             // 发出跳转命令
        #20;                       // 只需要维持一个周期
        jump_flag = 0;             // 恢复
        #60;                       // 看看是不是从 80001004 继续跑

        // --- 结束仿真 ---
        $stop;
    end

endmodule