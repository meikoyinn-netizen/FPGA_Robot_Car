`timescale 1ns / 1ps

// Synthesizable stub for Xilinx ILA IP.
// Replace with the real ILA IP by adding it to the Vivado project.
module ila_0 (
    input  wire        clk,
    input  wire [15:0] probe0,
    input  wire        probe1,
    input  wire        probe2,
    input  wire [31:0] probe3,
    input  wire [3:0]  probe4,
    input  wire        probe5,
    input  wire        probe6,
    input  wire [4:0]  probe7,
    input  wire        probe8
);
endmodule